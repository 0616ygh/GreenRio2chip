`ifndef _HEHE_CFG_VH_
`define _HEHE_CFG_VH_

// `define SYNTHESIS
// `define DPRAM64_2R1W
`ifndef SYNTHESIS
    // `define LSU_DEBUG
`endif // SYNTHESIS

`define LSU_V1

`endif // _HEHE_CFG_VH_
