`ifndef __UOP_ENCODING_PKG_SV__
`define __UOP_ENCODING_PKG_SV__

package uop_encoding_pkg;

   


endpackage

`endif